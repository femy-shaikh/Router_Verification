/************************************************************************
  
Copyright 2019 - Maven Silicon Softech Pvt Ltd.  
  
www.maven-silicon.com 
  
All Rights Reserved. 
This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd. 
It is not to be shared with or used by any third parties who have not enrolled for our paid 
training courses or received any written authorization from Maven Silicon.
  
Filename				:   router_wr_sequencer.sv

Description			:		Write sequencer class for Router 1x3
  
Author Name			:   Shanthi V A

Support e-mail	: 	For any queries, reach out to us on "techsupport_vm@maven-silicon.com" 

Version					:		1.0

************************************************************************/
class router_wr_sequencer extends uvm_sequencer #(write_xtn);

   // Factory registration using `uvm_component_utils
	 `uvm_component_utils(router_wr_sequencer)


   // Standard UVM Methods:
	 extern function new(string name = "router_wr_sequencer",uvm_component parent);
endclass

//-----------------  constructor new method  -------------------//
function router_wr_sequencer::new(string name="router_wr_sequencer",uvm_component parent);
	 super.new(name,parent);
endfunction

 

